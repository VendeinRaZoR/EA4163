module vmeout(
input R_
output [15:0] DOUT
);


endmodule 